library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity soc is
end soc;

architecture Behavioral of soc is

begin


end Behavioral;

